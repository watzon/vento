module main

import os

pub struct InputFile {
pub mut:
	filename string
	content_type string
	data string
}
